--top level vhdl
use library;
use conveyor;

1_conveyor:
	component conveyor
	generic map ();
	port map();
