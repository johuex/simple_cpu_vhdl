-- template for 1 of 10 conveyor
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

component conveyor is
generic ();
port ();
end component conveyor;